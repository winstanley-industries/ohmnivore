* Pulse Through RC Filter
* A 1kHz square wave (0-5V) drives an RC low-pass filter.
* The output shows the capacitor charging and discharging,
* rounding the square wave into a smoother waveform.

V1 in 0 PULSE(0 5 0 1n 1n 0.5m 1m)
R1 in out 1k
C1 out 0 1u

.TRAN 10u 3m 0 UIC
.PRINT TRAN V(in) V(out)
.END
