* Current Source with Resistor
I1 0 1 DC 0.001
R1 1 0 1k
.DC
.END
